* K544UD2A OPERATIONAL AMPLIFIER "MACROMODEL" SUBCIRCUIT
* VERSION 94/53dB@20kHz
* (REV N/A)      SUPPLY VOLTAGE: +/-15V
* CONNECTIONS:   NON-INVERTING INPUT
*                | INVERTING INPUT
*                | | POSITIVE POWER SUPPLY
*                | | | NEGATIVE POWER SUPPLY
*                | | | | OUTPUT
*                | | | | | FCORRECTION PIN 1
*                | | | | | | FCORRECTION PIN 8
*                | | | | | | |
.SUBCKT K544UD2A   In+ In- V+ V- OUT FC1 FC8
Cp1 OUT V- 3p
Cp2  FC1 V- 3p
Cp3 FC8 V-  3p 
Q2 N005 N001 V+ 0 PN
Q3 N001 N001 V+ 0 PN
Q12 N001 N001 V+ 0 PN
Q17 N006 N001 V+ 0 PN
Q4 N012 N005 N001 0 PN
Q13 N013 N006 N001 0 PN
Q5 N016 N015 N012 0 PN
Q14 N017 N015 N013 0 PN
Q8 N010 N010 N015 0 NP
J1 N005 In- N021 NJ
J18 N006 In+ N021 NJ
Q15 N017 N027 N035 0 NP
Q16 N035 N034 N042 0 NP
Q9 N024 N016 N027 0 NP
Q6 N016 N027 N034 0 NP
Q7 N034 N034 N041 0 NP
Q10 N031 N031 N040 0 NP
Q11 N040 N040 V- 0 NP
Q20 N037 N036 N044 0 NP
Q19 N021 N029 N037 0 NP
Q21 N021 N026 N029 0 NP
Q24 N026 N029 N036 0 NP
Q25 N036 N036 N045 0 NP
Q23 N023 N014 N026 0 NP
R1 N044 V- 230
R2 N045 V- 430
R3 N014 N023 110
R4 N010 N006 750
R5 N005 N010 750
R6 N009 N005 4k
R7 N027 N031 30k
R8 N042 V- 240
R9 N041 V- 240
Q26 N008 N002 V+ 0 PN
Q22 N014 N008 N002 0 PN
Q27 N008 N008 N015 0 NP
R10 V+ N002 1k6
R11 N006 N007 1k
R12 FC1 N006 200
Q28 N019 N023 N026 0 NP
R13 N015 N019 27k
R14 V+ N003 40k
D1 FC8 N003 DX
R15 FC8 N011 40k
D2 N015 N011 DX
C1 FC8 N017 12p 
J34 V+ N017 N018 NJ
Q38 V+ N018 N020 0 NP 
Q33 N007 N004 V+ 0 PN
R16 V+ N004 36
R19 N043 V- 36
Q41 N004 N020 N022 0 NP
R20 N022 OUT 36
R21 OUT N028 36
Q42 N043 N030 N028 0 PN
Q39 N020 N020 N025 0 NP
Q35 N020 N025 N030 0 NP
R17 N025 N030 40k
Q40 N036 N043 V- 0 NP
Q37 N039 N036 N047 0 NP
R18 N047 V- 240
Q31 N038 N036 N046 0 NP
R22 N046 V- 560
Q29 N032 N032 N036 0 NP
R23 N029 N032 6k6
Q30 N018 N029 N038 0 NP
Q36 N030 N033 N039 0 NP
Q32 V- N036 N033 0 PN 
R24 N019 N033 18k
D3 N017 N024 DX
* 3 (IN+)
* 2 (IN-)
* 1 (NC/FC)
* 8 (FC)
* 5 (NC)
.model NJ NJF Is=15p Beta=3.6m Vto=-1.5 cgs=3pF cgd=3pF lambda=10m kf=1e-16 af=0.3
.model NP NPN(BF=150 Cje=.25p Cjc=0.3p  VAF=100 tf=0.01n cjs=3p mjs=0.5 VTF=5 nf=1.0 )
.model PN LPNP(BF=35 Cje=.25p Cjc=1.p  VAF=50 tf=0.3n cjs=5.0p mjs=0.5 VTF=5 )
.model DX D(Is=2.52n Rs=.568 N=1.752 Cjo=0.4p M=.4 Tt=20n)
.ends K544UD2A

